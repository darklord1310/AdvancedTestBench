library verilog;
use verilog.vl_types.all;
entity adder_tb is
    generic(
        n               : integer := 4
    );
end adder_tb;
